*** SPICE deck for cell flop3{sch} from library cmoscells
*** Created on 星期五 六月 28, 2024 23:05:05
*** Last revised on 星期五 六月 28, 2024 23:14:40
*** Written on 星期五 六月 28, 2024 23:14:52 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: flop3{sch}
Mnmos@0 d clk net@6 gnd NMOS L=0.6U W=1.8U
Mnmos@1 net@6 net@8 gnd gnd NMOS L=0.6U W=1.8U
Mnmos@2 net@11 clk gnd gnd NMOS L=0.6U W=1.8U
Mnmos@3 d net@11 net@38 gnd NMOS L=0.6U W=1.8U
Mnmos@4 net@38 net@31 gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 net@7 net@11 d vdd PMOS L=0.6U W=3.6U
Mpmos@1 vdd net@8 net@7 vdd PMOS L=0.6U W=3.6U
Mpmos@2 vdd clk net@11 vdd PMOS L=0.6U W=3.6U
Mpmos@3 net@39 clk d vdd PMOS L=0.6U W=3.6U
Mpmos@4 vdd net@31 net@39 vdd PMOS L=0.6U W=3.6U

* Spice Code nodes in cell cell 'flop3{sch}'
vdd vdd 0 DC 5
va clk 0 PULSE(0 5 0n 1n 1n 20n 40n)
vb d 0 DC pwl 30n 0 31n 5 105n 5 106n 0
.tran 200n
.include c5_models.txt
.END
