*** SPICE deck for cell MUX{lay} from library cmoscells
*** Created on 星期五 六月 28, 2024 21:31:59
*** Last revised on 星期六 六月 29, 2024 22:27:02
*** Written on 星期六 六月 29, 2024 22:27:09 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: MUX{lay}
Mnmos@0 net@1 C gnd gnd NMOS L=0.6U W=1.8U AS=30.24P AD=4.86P PS=46.2U PD=9U
Mnmos@1 B net@1 Q gnd NMOS L=0.6U W=1.8U AS=4.86P AD=4.86P PS=9U PD=9U
Mnmos@2 Q C A gnd NMOS L=0.6U W=1.8U AS=4.86P AD=4.86P PS=9U PD=9U
Mpmos@0 net@1 C vdd vdd PMOS L=0.6U W=3.6U AS=38.88P AD=4.86P PS=50.4U PD=9U
Mpmos@1 B C Q vdd PMOS L=0.6U W=3.6U AS=4.86P AD=4.86P PS=9U PD=9U
Mpmos@2 Q net@1 A vdd PMOS L=0.6U W=3.6U AS=4.86P AD=4.86P PS=9U PD=9U

* Spice Code nodes in cell cell 'MUX{lay}'
vdd vdd 0 DC 5
va A 0 PULSE(0 5 0n 1n 1n 20n 40n)
vb B 0 DC pwl 30n 0 31n 5 55n 5 56n 0 80n 0 81n 5 115n 5 116n 0
vc c 0 DC pwl 25n 0 26n 5 105n 5 106n 0
.tran 200n
.include C5_models.txt
.END
