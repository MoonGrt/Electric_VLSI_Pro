*** SPICE deck for cell flop{sch} from library blood_oxygen
*** Created on 星期三 十二月 20, 2000 00:40:01
*** Last revised on 星期五 六月 28, 2024 10:47:58
*** Written on 星期五 六月 28, 2024 10:48:02 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: blood_oxygen:flop{sch}
Mnmos@0 gnd net@2 net@32 gnd SPICE-Model L=0.6U W=1.8U
Mnmos@1 net@10 ph2b net@32 gnd N L=0.6U W=1.8U
Mnmos@2 net@2 net@10 gnd gnd N L=0.6U W=1.8U
Mnmos@3 net@10 ph2 d gnd NMOS L=0.6U W=1.8U
Mnmos@4 gnd net@53 net@62 gnd N L=0.6U W=1.8U
Mnmos@5 net@14 ph1b net@62 gnd N L=0.6U W=1.8U
Mnmos@6 net@53 net@14 gnd gnd N L=0.6U W=1.8U
Mnmos@7 q net@14 gnd gnd N L=0.6U W=1.8U
Mnmos@8 net@14 ph1 net@2 gnd N L=0.6U W=1.8U
Mpmos@0 net@43 ph2 net@10 vdd P L=0.6U W=3.6U
Mpmos@1 net@43 net@2 vdd vdd P L=0.6U W=3.6U
Mpmos@2 vdd net@10 net@2 vdd P L=0.6U W=3.6U
Mpmos@3 d ph2b net@10 vdd PMOS L=0.6U W=3.6U
Mpmos@4 net@12 ph1 net@14 vdd P L=0.6U W=3.6U
Mpmos@5 net@12 net@53 vdd vdd P L=0.6U W=3.6U
Mpmos@6 vdd net@14 net@53 vdd P L=0.6U W=3.6U
Mpmos@7 vdd net@14 q vdd P L=0.6U W=3.6U
Mpmos@8 net@2 ph1b net@14 vdd P L=0.6U W=3.6U
.END
