*** SPICE deck for cell MUX_sim{lay} from library cmoscells
*** Created on 星期一 七月 01, 2024 06:53:54
*** Last revised on 星期一 七月 01, 2024 06:57:24
*** Written on 星期一 七月 01, 2024 07:26:47 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__MUX FROM CELL MUX{lay}
.SUBCKT cmoscells__MUX A B C gnd Q vdd
Mnmos@0 net@3 C gnd gnd NMOS L=0.4U W=1.2U AS=13.44P AD=2.16P PS=30.8U PD=6U
Mnmos@1 B net@3 Q gnd NMOS L=0.4U W=1.2U AS=2.16P AD=2.16P PS=6U PD=6U
Mnmos@2 Q C A gnd NMOS L=0.4U W=1.2U AS=2.16P AD=2.16P PS=6U PD=6U
Mpmos@0 net@3 C vdd vdd PMOS L=0.4U W=2.4U AS=17.28P AD=2.16P PS=33.6U PD=6U
Mpmos@1 B C Q vdd PMOS L=0.4U W=2.4U AS=2.16P AD=2.16P PS=6U PD=6U
Mpmos@2 Q net@3 A vdd PMOS L=0.4U W=2.4U AS=2.16P AD=2.16P PS=6U PD=6U
.ENDS cmoscells__MUX

*** TOP LEVEL CELL: MUX_sim{lay}
XMUX@0 A B C gnd Q vdd cmoscells__MUX

* Spice Code nodes in cell cell 'MUX_sim{lay}'
vdd vdd 0 DC 5
va A 0 PULSE(0 5 0n 1n 1n 20n 40n)
vb B 0 DC pwl 30n 0 31n 5 55n 5 56n 0 80n 0 81n 5 115n 5 116n 0
vc c 0 DC pwl 25n 0 26n 5 105n 5 106n 0
.tran 200n
.include C5_models.txt
.END
