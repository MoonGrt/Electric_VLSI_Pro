*** SPICE deck for cell INV_sim{lay} from library cmoscells
*** Created on 星期一 七月 01, 2024 06:53:01
*** Last revised on 星期一 七月 01, 2024 07:00:23
*** Written on 星期一 七月 01, 2024 07:24:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__INV FROM CELL INV{lay}
.SUBCKT cmoscells__INV gnd in out vdd
Mnmos@0 out in gnd gnd NMOS L=0.4U W=1.2U AS=2.32P AD=1.98P PS=8.6U PD=5.8U
Mpmos@0 out in vdd vdd PMOS L=0.4U W=2.4U AS=3.64P AD=1.98P PS=11U PD=5.8U
.ENDS cmoscells__INV

*** TOP LEVEL CELL: INV_sim{lay}
XINV@0 gnd in out vdd cmoscells__INV

* Spice Code nodes in cell cell 'INV_sim{lay}'
vdd vdd 0 DC 5
va in 0 PULSE(0 5 0n 1n 1n 20n 40n)
.tran 200n
.include C5_models.txt
.END
