*** SPICE deck for cell std_inv{sch} from library blood_oxygen
*** Created on 星期二 十二月 19, 2000 08:56:10
*** Last revised on 星期五 六月 28, 2024 10:52:19
*** Written on 星期五 六月 28, 2024 10:52:22 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: blood_oxygen:std_inv{sch}
Mnmos@0 y a gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd a y vdd PMOS L=0.6U W=3.6U

* Spice Code nodes in cell cell 'blood_oxygen:std_inv{sch}'
vdd vdd 0 DC 5
vin a 0 DC pwl 10ns 0 20ns 5 50ns 5 60ns 0
cload y 0 250fF
.measure tran tf trig v(out) val=4.5 fall=1 td=8ns targ v(out) val=0.5 fall=1
.measure tran tr trig v(out) val=0.5 rise=1 td=50ns targ v(out) val=4.5 rise=1
.tran 0 0.1us
.include F:\Study\DIC\Lab\Lab2\Lab2_files\C5_models.txt
.END
