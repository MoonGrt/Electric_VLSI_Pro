*** SPICE deck for cell NAND{lay} from library blood_oxygen
*** Created on 星期四 六月 27, 2024 16:43:57
*** Last revised on 星期四 六月 27, 2024 17:08:45
*** Written on 星期四 六月 27, 2024 17:08:51 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND{lay}
Mnmos@0 gnd B net@20 gnd NMOS L=2U W=10U AS=30P AD=250P PS=16U PD=115U
Mnmos@1 net@20 A AB gnd N L=2U W=10U AS=58.333P AD=30P PS=25U PD=16U
Mpmos@0 vdd B AB vdd PMOS L=2U W=10U AS=58.333P AD=162.5P PS=25U PD=75U
Mpmos@1 AB A vdd vdd PMOS L=2U W=10U AS=162.5P AD=58.333P PS=75U PD=25U
.END
