*** SPICE deck for cell add1{sch} from library cmoscells
*** Created on 星期五 六月 28, 2024 23:16:38
*** Last revised on 星期六 六月 29, 2024 18:18:10
*** Written on 星期日 六月 30, 2024 20:12:24 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__std_inv FROM CELL std_inv{sch}
.SUBCKT cmoscells__std_inv a y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 y a gnd gnd NMOS L=0.4U W=1.2U
Mpmos@0 vdd a y vdd PMOS L=0.4U W=2.4U
.ENDS cmoscells__std_inv

.global gnd vdd

*** TOP LEVEL CELL: add1{sch}
Mnmos@7 net@87 gnd net@73 gnd NMOS L=0.4U W=1.2U
Mnmos@9 net@82 A net@87 gnd NMOS L=0.4U W=1.2U
Mnmos@10 net@82 C net@70 gnd NMOS L=0.4U W=1.2U
Mnmos@11 net@70 A net@73 gnd NMOS L=0.4U W=1.2U
Mnmos@15 net@70 gnd net@73 gnd NMOS L=0.4U W=1.2U
Mnmos@16 net@241 C gnd gnd NMOS L=0.4U W=1.2U
Mnmos@17 net@241 A gnd gnd NMOS L=0.4U W=1.2U
Mnmos@18 net@241 gnd gnd gnd NMOS L=0.4U W=1.2U
Mnmos@19 net@116 net@82 net@241 gnd NMOS L=0.4U W=1.2U
Mnmos@20 net@116 C net@247 gnd NMOS L=0.4U W=1.2U
Mnmos@21 net@247 A net@249 gnd NMOS L=0.4U W=1.2U
Mnmos@22 net@249 gnd gnd gnd NMOS L=0.4U W=1.2U
Mpmos@10 vdd C net@104 vdd PMOS L=0.4U W=2.4U
Mpmos@11 vdd A net@104 vdd PMOS L=0.4U W=2.4U
Mpmos@12 vdd gnd net@104 vdd PMOS L=0.4U W=2.4U
Mpmos@13 net@104 net@82 net@116 vdd PMOS L=0.4U W=2.4U
Mpmos@14 net@104 C net@107 vdd PMOS L=0.4U W=2.4U
Mpmos@15 net@107 A net@108 vdd PMOS L=0.4U W=2.4U
Mpmos@16 net@108 gnd net@116 vdd PMOS L=0.4U W=2.4U
Mpmos@17 vdd A net@200 vdd PMOS L=0.4U W=2.4U
Mpmos@18 net@200 A net@195 vdd PMOS L=0.4U W=2.4U
Mpmos@19 net@195 gnd net@82 vdd PMOS L=0.4U W=2.4U
Mpmos@20 vdd gnd net@200 vdd PMOS L=0.4U W=2.4U
Mpmos@21 net@200 C net@82 vdd PMOS L=0.4U W=2.4U
Xstd_inv@0 net@82 C1 cmoscells__std_inv
Xstd_inv@1 net@116 S cmoscells__std_inv

* Spice Code nodes in cell cell 'add1{sch}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 11n 5 50n 5 51n 0 90n 0 91n 5 130n 5 131n 0 170n 0 171n 5
vb B 0 DC 5
vc C 0 DC pwl 30n 0 31n 5 105n 5 106n 0
.tran 200n
.include c5_models.txt
.END
