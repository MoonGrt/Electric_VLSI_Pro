*** SPICE deck for cell add1_sim{lay} from library cmoscells
*** Created on 星期一 七月 01, 2024 07:07:57
*** Last revised on 星期一 七月 01, 2024 07:11:04
*** Written on 星期一 七月 01, 2024 07:33:45 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__add1 FROM CELL add1{lay}
.SUBCKT cmoscells__add1 A B C C1 gnd S vdd
Mnmos@0 gnd B net@134 gnd NMOS L=0.4U W=1.2U AS=1.52P AD=7.469P PS=4.133U PD=16.743U
Mnmos@1 net@134 A gnd gnd NMOS L=0.4U W=1.2U AS=7.469P AD=1.52P PS=16.743U PD=4.133U
Mnmos@2 net@83 C net@134 gnd NMOS L=0.4U W=1.2U AS=1.52P AD=2.58P PS=4.133U PD=5.7U
Mnmos@4 C1 net@83 gnd gnd NMOS L=0.4U W=1.2U AS=7.469P AD=2.16P PS=16.743U PD=6U
Mnmos@6 net@253 B net@83 gnd NMOS L=0.4U W=1.2U AS=2.58P AD=0.72P PS=5.7U PD=2.4U
Mnmos@7 gnd A net@253 gnd NMOS L=0.4U W=1.2U AS=0.72P AD=7.469P PS=2.4U PD=16.743U
Mnmos@13 net@209 A net@285 gnd NMOS L=0.4U W=1.2U AS=0.72P AD=1.824P PS=2.4U PD=4.32U
Mnmos@14 net@273 A net@209 gnd NMOS L=0.4U W=1.2U AS=1.824P AD=1.32P PS=4.32U PD=3.4U
Mnmos@15 net@209 B net@273 gnd NMOS L=0.4U W=1.2U AS=1.32P AD=1.824P PS=3.4U PD=4.32U
Mnmos@17 gnd net@83 net@273 gnd NMOS L=0.4U W=1.2U AS=1.32P AD=7.469P PS=3.4U PD=16.743U
Mnmos@18 net@273 C net@209 gnd NMOS L=0.4U W=1.2U AS=1.824P AD=1.32P PS=4.32U PD=3.4U
Mnmos@19 net@285 B net@286 gnd NMOS L=0.4U W=1.2U AS=0.72P AD=0.72P PS=2.4U PD=2.4U
Mnmos@20 net@286 C gnd gnd NMOS L=0.4U W=1.2U AS=7.469P AD=0.72P PS=16.743U PD=2.4U
Mnmos@21 S net@209 gnd gnd NMOS L=0.4U W=1.2U AS=7.469P AD=2.16P PS=16.743U PD=6U
Mpmos@0 net@85 A vdd vdd PMOS L=0.4U W=2.4U AS=9.909P AD=2.64P PS=17.886U PD=4.6U
Mpmos@2 net@84 A net@83 vdd PMOS L=0.4U W=2.4U AS=2.58P AD=1.44P PS=5.7U PD=3.6U
Mpmos@3 net@85 B net@84 vdd PMOS L=0.4U W=2.4U AS=1.44P AD=2.64P PS=3.6U PD=4.6U
Mpmos@4 vdd B net@85 vdd PMOS L=0.4U W=2.4U AS=2.64P AD=9.909P PS=4.6U PD=17.886U
Mpmos@9 net@83 net@179 net@85 vdd PMOS L=0.4U W=2.4U AS=2.64P AD=2.58P PS=4.6U PD=5.7U
Mpmos@10 C1 net@83 vdd vdd PMOS L=0.4U W=2.4U AS=9.909P AD=2.16P PS=17.886U PD=6U
Mpmos@11 net@210 net@83 net@209 vdd PMOS L=0.4U W=2.4U AS=1.824P AD=2.88P PS=4.32U PD=5.28U
Mpmos@13 net@210 B vdd vdd PMOS L=0.4U W=2.4U AS=9.909P AD=2.88P PS=17.886U PD=5.28U
Mpmos@14 vdd A net@210 vdd PMOS L=0.4U W=2.4U AS=2.88P AD=9.909P PS=5.28U PD=17.886U
Mpmos@15 vdd C net@210 vdd PMOS L=0.4U W=2.4U AS=2.88P AD=9.909P PS=5.28U PD=17.886U
Mpmos@16 net@225 A net@210 vdd PMOS L=0.4U W=2.4U AS=2.88P AD=1.44P PS=5.28U PD=3.6U
Mpmos@17 net@226 B net@225 vdd PMOS L=0.4U W=2.4U AS=1.44P AD=1.44P PS=3.6U PD=3.6U
Mpmos@18 net@227 C net@226 vdd PMOS L=0.4U W=2.4U AS=1.44P AD=3.84P PS=3.6U PD=8U
Mpmos@19 S net@209 vdd vdd PMOS L=0.4U W=2.4U AS=9.909P AD=2.16P PS=17.886U PD=6U
.ENDS cmoscells__add1

*** TOP LEVEL CELL: add1_sim{lay}
Xadd1@1 A B C C1 gnd S vdd cmoscells__add1

* Spice Code nodes in cell cell 'add1_sim{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 11n 5 50n 5 51n 0 90n 0 91n 5 130n 5 131n 0 170n 0 171n 5
vb B 0 DC 5
vc C 0 DC pwl 30n 0 31n 5 105n 5 106n 0
.tran 200n
.include c5_models.txt
.END
