*** SPICE deck for cell INV_sim{sch} from library cmoscells
*** Created on 星期一 七月 01, 2024 06:52:37
*** Last revised on 星期一 七月 01, 2024 06:58:48
*** Written on 星期一 七月 01, 2024 15:07:53 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__INV FROM CELL INV{sch}
.SUBCKT cmoscells__INV in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=0.6U W=1.8U
Mpmos@0 vdd in out vdd PMOS L=0.6U W=3.6U
.ENDS cmoscells__INV

.global gnd vdd

*** TOP LEVEL CELL: INV_sim{sch}
XINV@0 in out cmoscells__INV

* Spice Code nodes in cell cell 'INV_sim{sch}'
vdd vdd 0 DC 5
va in 0 PULSE(0 5 0n 1n 1n 20n 40n)
.tran 200n
.include C5_models.txt
.END
