*** SPICE deck for cell XOR_sim{lay} from library cmoscells
*** Created on 星期一 七月 01, 2024 07:05:00
*** Last revised on 星期一 七月 01, 2024 07:32:05
*** Written on 星期一 七月 01, 2024 07:32:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__XOR FROM CELL XOR{lay}
.SUBCKT cmoscells__XOR A B gnd vdd XOR
Mnmos@0 net@86 A XOR gnd NMOS L=0.4U W=2U AS=2.2P AD=2.7P PS=4.2U PD=5.7U
Mnmos@3 gnd B net@86 gnd NMOS L=0.4U W=2U AS=2.7P AD=7.95P PS=5.7U PD=16.7U
Mnmos@4 gnd A net@94 gnd NMOS L=0.4U W=2U AS=3.2P AD=7.95P PS=7.2U PD=16.7U
Mnmos@5 net@45 B gnd gnd NMOS L=0.4U W=2U AS=7.95P AD=3.2P PS=16.7U PD=7.2U
Mnmos@6 net@86 net@94 gnd gnd NMOS L=0.4U W=2U AS=7.95P AD=2.7P PS=16.7U PD=5.7U
Mnmos@7 XOR net@45 net@86 gnd NMOS L=0.4U W=2U AS=2.7P AD=2.2P PS=5.7U PD=4.2U
Mpmos@1 net@98 net@45 XOR vdd PMOS L=0.4U W=2U AS=2.2P AD=1.2P PS=4.2U PD=3.2U
Mpmos@5 net@45 B vdd vdd PMOS L=0.4U W=2U AS=8.45P AD=3.2P PS=18.2U PD=7.2U
Mpmos@6 vdd A net@98 vdd PMOS L=0.4U W=2U AS=1.2P AD=8.45P PS=3.2U PD=18.2U
Mpmos@7 vdd A net@94 vdd PMOS L=0.4U W=2U AS=3.2P AD=8.45P PS=7.2U PD=18.2U
Mpmos@9 XOR net@94 net@154 vdd PMOS L=0.4U W=2U AS=1.2P AD=2.2P PS=3.2U PD=4.2U
Mpmos@10 net@154 B vdd vdd PMOS L=0.4U W=2U AS=8.45P AD=1.2P PS=18.2U PD=3.2U
.ENDS cmoscells__XOR

*** TOP LEVEL CELL: XOR_sim{lay}
XXOR@0 A B gnd vdd XOR cmoscells__XOR

* Spice Code nodes in cell cell 'XOR_sim{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 0 5 100n 5 110n 0
.tran 200n
.include c5_models.txt
.END
