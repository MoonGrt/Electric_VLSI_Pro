*** SPICE deck for cell NAND_sim{sch} from library cmoscells
*** Created on 星期六 一月 16, 2010 05:31:02
*** Last revised on 星期四 六月 27, 2024 16:35:44
*** Written on 星期五 六月 28, 2024 22:35:56 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__NAND FROM CELL NAND{sch}
.SUBCKT cmoscells__NAND A AB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AB A net@20 gnd NMOS L=0.6U W=3U
Mnmos@1 AB A vdd vdd PMOS L=0.6U W=3U
Mnmos@2 net@20 B gnd gnd NMOS L=0.6U W=3U
Mpmos@0 AB B vdd vdd PMOS L=0.6U W=3U
.ENDS cmoscells__NAND

.global gnd vdd

*** TOP LEVEL CELL: NAND_sim{sch}
XNAND@0 A AB B cmoscells__NAND

* Spice Code nodes in cell cell 'NAND_sim{sch}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.measure tran tf trig v(AB) val=4.5 fall=1 td=4ns targ v(AB) val=0.5 fall=1
.measure tran tr trig v(AB) val=0.5 rise=1 td=4ns targ v(AB) val=4.5 rise=1
.tran 200n
.include C5_models.txt
.END
