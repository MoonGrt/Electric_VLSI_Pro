*** SPICE deck for cell NAND_sim{lay} from library cmoscells
*** Created on 星期四 六月 27, 2024 16:19:20
*** Last revised on 星期四 六月 27, 2024 21:09:46
*** Written on 星期一 七月 01, 2024 07:28:45 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT cmoscells__NAND FROM CELL NAND{lay}
.SUBCKT cmoscells__NAND A AB B gnd vdd
Mnmos@0 gnd B net@20 gnd NMOS L=0.4U W=2U AS=1.2P AD=10P PS=3.2U PD=23U
Mnmos@1 net@20 A AB gnd NMOS L=0.4U W=2U AS=2.333P AD=1.2P PS=5U PD=3.2U
Mpmos@0 vdd B AB vdd PMOS L=0.4U W=2U AS=2.333P AD=6.5P PS=5U PD=15U
Mpmos@1 AB A vdd vdd PMOS L=0.4U W=2U AS=6.5P AD=2.333P PS=15U PD=5U
.ENDS cmoscells__NAND

*** TOP LEVEL CELL: NAND_sim{lay}
XNAND@2 A AB B gnd vdd cmoscells__NAND

* Spice Code nodes in cell cell 'NAND_sim{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.measure tran tf trig v(AB) val=4.5 fall=1 td=4ns targ v(AB) val=0.5 fall=1
.measure tran tr trig v(AB) val=0.5 rise=1 td=4ns targ v(AB) val=4.5 rise=1
.tran 200n
.include C5_models.txt
.END
